`timescale 1ns / 1ps

module Signal_Classifier (
    input wire clk,         // 100kHz �ý��� Ŭ��
    input wire rst_n,       // Reset
    input wire btn_in,      // Debounced Button Input (H: Pressed)
    
    output reg valid,       // 1: �ǵ� �Ϸ� (��ư �� �� 1Ŭ�� Pulse)
    output reg is_long      // 0: Short, 1: Long (valid�� ���� ��ȿ)
);

    // =========================================================================
    // 1. �Ķ���� ���� (100kHz ����)
    // =========================================================================
    // Long Press �Ǵ� ����: 300ms
    // 100,000Hz * 0.3s = 30,000 Ticks
    parameter LONG_PRESS_TH = 30000; 

    // =========================================================================
    // 2. ���� ����
    // =========================================================================
    reg [31:0] press_cnt;
    reg btn_prev; // Edge �����

    // =========================================================================
    // 3. ���� ����
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            press_cnt <= 0;
            btn_prev <= 0;
            valid <= 0;
            is_long <= 0;
        end else begin
            valid <= 0; // Pulse �ʱ�ȭ
            btn_prev <= btn_in;

            if (btn_in == 1'b1) begin
                // A. ��ư ������ ��: �ð� ����
                // Overflow �����ϸ� ī����
                if (press_cnt < LONG_PRESS_TH + 10) 
                    press_cnt <= press_cnt + 1;
            end 
            else begin
                // B. ��ư�� ���� �� (Falling Edge)
                if (btn_prev == 1'b1) begin
                    valid <= 1'b1; // ��� ���Դٰ� �˸�
                    
                    // C. �ð� �Ǻ�
                    if (press_cnt >= LONG_PRESS_TH) is_long <= 1'b1;
                    else                            is_long <= 1'b0;
                end
                
                // ī���� �ʱ�ȭ
                press_cnt <= 0;
            end
        end
    end

endmodule