`timescale 1ns / 1ps

module tb_Button_Debouncer;

    // =========================================================================
    // 1. ���� �� DUT ����
    // =========================================================================
    reg clk;
    reg rst_n;
    reg btn_in;
    wire btn_out;

    // 100kHz ȯ�� ����
    parameter TEST_CLK_FREQ = 100_000;
    parameter TEST_DEBOUNCE_MS = 20;

    Button_Debouncer #(
        .CLK_FREQ(TEST_CLK_FREQ), 
        .DEBOUNCE_MS(TEST_DEBOUNCE_MS)
    ) uut (
        .clk(clk),
        .rst_n(rst_n),
        .btn_in(btn_in),
        .btn_out(btn_out)
    );

    // =========================================================================
    // 2. 100kHz Ŭ�� ���� (Divider ���� ���� ����)
    // =========================================================================
    initial begin
        clk = 0;
    end
    
    // 5000ns(5us)���� ���� -> �ֱ� 10us -> 100kHz
    always #5000 clk = ~clk; 

    // =========================================================================
    // 3. �׽�Ʈ �ó�����
    // =========================================================================
    initial begin
        $display("=== Simulation Start (100kHz Clock) ===");
        
        // �ʱ�ȭ
        rst_n = 0;
        btn_in = 0;
        #2_000_000; // 2ms ���
        rst_n = 1;
        #2_000_000;

        // ---------------------------------------------------------------------
        // Case 1: ª�� ������ (5ms) -> ���õǾ�� ��
        // ---------------------------------------------------------------------
        $display("[Time: %t] Noise Injection (5ms)", $time);
        btn_in = 1; 
        #5_000_000; // 5ms ���� (������ 20ms �̸�)
        btn_in = 0;
        
        #30_000_000; // ����� ��� (30ms)

        if (btn_out == 0) $display(" -> PASS: Noise Ignored");
        else              $display(" -> FAIL: Noise Detected");

        // ---------------------------------------------------------------------
        // Case 2: ���� �Է� (30ms) -> �νĵǾ�� ��
        // ---------------------------------------------------------------------
        $display("[Time: %t] Stable Press (30ms)", $time);
        btn_in = 1;
        #30_000_000; // 30ms ���� (������ 20ms �̻�)
        
        if (btn_out == 1) $display(" -> PASS: Signal Detected");
        else              $display(" -> FAIL: Signal Missed");

        // ---------------------------------------------------------------------
        // Case 3: ��ư �� -> ���� Ȯ��
        // ---------------------------------------------------------------------
        btn_in = 0;
        #30_000_000;
        
        if (btn_out == 0) $display(" -> PASS: Release Detected");
        else              $display(" -> FAIL: Release Failed");

        $display("=== Simulation End ===");
        $finish;
    end

endmodule