`timescale 1ns / 1ps

module tb_top;

    // Inputs
    reg clk;
    reg rst_n;
    reg [3:0] key_val;
    reg key_trig;

    // Outputs
    wire lcd_rs;
    wire lcd_rw;
    wire lcd_e;
    wire [7:0] lcd_data;
    wire piezo_out;  // [����] Top.v�� ��Ʈ��� ��ġ��Ŵ
    wire [3:0] led;

    // Instantiate the Unit Under Test (UUT)
    Top uut (
        .clk(clk), 
        .rst_n(rst_n), 
        .key_val(key_val), 
        .key_trig(key_trig), 
        .lcd_rs(lcd_rs), 
        .lcd_rw(lcd_rw), 
        .lcd_e(lcd_e), 
        .lcd_data(lcd_data), 
        .piezo_out(piezo_out), // [����] ���� �߻��ϴ� �κ� �ذ�
        .led(led)
    );

    // Clock Generation (100MHz)
    always #5 clk = ~clk;

    initial begin
        // Initialize Inputs
        clk = 0;
        rst_n = 0;
        key_val = 0;
        key_trig = 0;

        // Wait 100 ns for global reset to finish
        #100;
        rst_n = 1;
        #100;
        
        // --- �׽�Ʈ �ó����� ���� ---
        
        // 1. ��(Dot) �Է� (A�� �պκ�)
        key_val = 4'd1; // KEY_DOT
        key_trig = 1;   // ��ư ����
        #20;
        key_trig = 0;   // ��ư ��
        #100000;        // ó�� ���

        // 2. ��(Dash) �Է� (A�� �޺κ�)
        key_val = 4'd2; // KEY_DASH
        key_trig = 1;
        #20;
        key_trig = 0;
        #100000;

        // 3. ��� (�ڵ� ���� Ʈ���� Ȯ��)
        #50000000; // ����� �ð� ���
        
        $stop;
    end
      
endmodule