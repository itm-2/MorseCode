module Top(
    input wire clk,
    input wire rst_n,
    
    // Ű�е� ��� ��� ���� �Է� ���� (����ġ 4��, ��ư 1�� ��)
    input wire [3:0] key_val,  // Ű �� (��: ����ġ)
    input wire key_trig,       // Ű �Է� ��ȣ (��: ��ư)
    
    output wire lcd_rs,
    output wire lcd_rw,
    output wire lcd_e,
    output wire [7:0] lcd_data,
    
    output wire piezo_out,     // ���� ���
    output wire [3:0] led      // LED ���
    );

    // --- UI ��� ���� ��ȣ ---
    wire ui_piezo_enable;
    wire [15:0] ui_freq;
    wire ui_req_mode_change;
    wire [3:0] ui_version;
    wire ui_is_error;
    wire [3:0] ui_led_out;

    // --- DecodeUI �ν��Ͻ� ---
    DecodeUI u_ui (
        .clk(clk),
        .rst_n(rst_n),
        .is_active(1'b1),        
        .key_valid(key_trig),    // ��ư ������ �Է� ��ȿ
        .k_data(key_val),        // ����ġ ���� �����ͷ� ���
        .key_pressed(key_trig),  // ��ư ���� ����
        
        // LCD
        .lcd_rs(lcd_rs),
        .lcd_rw(lcd_rw),
        .lcd_e(lcd_e),
        .lcd_data(lcd_data),
        
        // Sound & LED & Status (���� ���� ��Ʈ�� ���� �Ϸ�)
        .piezo(ui_piezo_enable), 
        .piezo_freq(ui_freq),    
        .req_mode_change(ui_req_mode_change),
        .ui_version(ui_version),
        .is_error(ui_is_error),  
        .led_out(ui_led_out)     
    );

    // --- LED ��� ---
    // ������ ��ü ����, �ƴϸ� UI���� �� �� ���
    assign led = ui_is_error ? 4'b1111 : ui_led_out;

    // --- �ǿ��� �Ҹ� �߻��� (Tone Generator) ---
    // UI���� ���� ���ļ�(ui_freq)�� �Ҹ� ���
    reg [31:0] tone_cnt;
    reg tone_clk;
    
    // 100MHz Ŭ�� ���� (���忡 �°� ���� ����)
    wire [31:0] toggle_value = (ui_freq > 0) ? (100_000_000 / ui_freq) / 2 : 32'd100000;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            tone_cnt <= 0;
            tone_clk <= 0;
        end else if (ui_piezo_enable) begin
            if (tone_cnt >= toggle_value) begin
                tone_cnt <= 0;
                tone_clk <= ~tone_clk;
            end else begin
                tone_cnt <= tone_cnt + 1;
            end
        end else begin
            tone_cnt <= 0;
            tone_clk <= 0;
        end
    end

    assign piezo_out = tone_clk;

endmodule