`timescale 1ns / 1ps

module ButtonMorseInput #(
    parameter DEBOUNCE_CYCLES = 250_000           // 10ms ��ٿ
)(
    input  wire        clk,
    input  wire        rst_n,
    input  wire [4:0]  btn,                        // btn[0]=��ư1, btn[1]=��ư2, btn[2]=PAUSE, btn[3]=CLEAR
    
    input wire [31:0] LONG_KEY_CYCLES,             // 500ms (DASH ����)
    input wire [31:0] DIT_GAP_CYCLES,              // 250ms (�ڵ� �ݺ� �ֱ�)
    
    output reg         key_valid,
    output reg  [10:0] key_packet,
    
    output reg         btn1_held,                  // ��ư1 ������ �� (�ǿ�����)
    output reg         btn2_dot_pulse              // ��ư2 DOT �޽� (�ǿ�����)
);

    localparam TYPE_KEY = 3'b001;
    localparam KEY_DOT   = 8'd1;
    localparam KEY_DASH  = 8'd2;
    localparam KEY_CLEAR = 8'd11;
    localparam KEY_PAUSE = 8'd12;

    //==========================================================================
    // 1. Synchronizer (2-stage flip-flop)
    //==========================================================================
    reg [1:0] b0_sync, b1_sync, b2_sync, b3_sync;
    
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            b0_sync <= 2'b00;
            b1_sync <= 2'b00;
            b2_sync <= 2'b00;
            b3_sync <= 2'b00;
        end else begin
            b0_sync <= {b0_sync[0], btn[0]};
            b1_sync <= {b1_sync[0], btn[1]};
            b2_sync <= {b2_sync[0], btn[2]};
            b3_sync <= {b3_sync[0], btn[3]};
        end
    end

    //==========================================================================
    // 2. Debouncer for btn[0] (��ư1)
    //==========================================================================
    reg        b0_stable;
    reg [31:0] b0_counter;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            b0_stable <= 1'b0;
            b0_counter <= 32'd0;
        end else begin
            if(b0_sync[1] != b0_stable) begin
                if(b0_counter >= DEBOUNCE_CYCLES) begin
                    b0_stable <= b0_sync[1];
                    b0_counter <= 32'd0;
                end else begin
                    b0_counter <= b0_counter + 1;
                end
            end else begin
                b0_counter <= 32'd0;
            end
        end
    end

    //==========================================================================
    // 3. Debouncer for btn[1] (��ư2)
    //==========================================================================
    reg        b1_stable;
    reg [31:0] b1_counter;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            b1_stable <= 1'b0;
            b1_counter <= 32'd0;
        end else begin
            if(b1_sync[1] != b1_stable) begin
                if(b1_counter >= DEBOUNCE_CYCLES) begin
                    b1_stable <= b1_sync[1];
                    b1_counter <= 32'd0;
                end else begin
                    b1_counter <= b1_counter + 1;
                end
            end else begin
                b1_counter <= 32'd0;
            end
        end
    end

    //==========================================================================
    // 4. Debouncer for btn[2] (PAUSE)
    //==========================================================================
    reg        b2_stable;
    reg [31:0] b2_counter;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            b2_stable <= 1'b0;
            b2_counter <= 32'd0;
        end else begin
            if(b2_sync[1] != b2_stable) begin
                if(b2_counter >= DEBOUNCE_CYCLES) begin
                    b2_stable <= b2_sync[1];
                    b2_counter <= 32'd0;
                end else begin
                    b2_counter <= b2_counter + 1;
                end
            end else begin
                b2_counter <= 32'd0;
            end
        end
    end

    //==========================================================================
    // 5. Debouncer for btn[3] (CLEAR)
    //==========================================================================
    reg        b3_stable;
    reg [31:0] b3_counter;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            b3_stable <= 1'b0;
            b3_counter <= 32'd0;
        end else begin
            if(b3_sync[1] != b3_stable) begin
                if(b3_counter >= DEBOUNCE_CYCLES) begin
                    b3_stable <= b3_sync[1];
                    b3_counter <= 32'd0;
                end else begin
                    b3_counter <= b3_counter + 1;
                end
            end else begin
                b3_counter <= 32'd0;
            end
        end
    end

    //==========================================================================
    // 6. ��ư ���� ����
    //==========================================================================
    reg        b0_prev;
    reg [31:0] b0_hold_counter;
    reg        b0_long_triggered;

    reg        b1_prev;
    reg [31:0] b1_repeat_counter;
    reg        b1_first_dot_sent;

    reg        b2_prev;
    reg        b3_prev;

    wire b0_pressed = (b0_stable && !b0_prev);
    wire b0_released = (!b0_stable && b0_prev);
    wire b0_holding = b0_stable;

    wire b1_pressed = (b1_stable && !b1_prev);
    wire b1_released = (!b1_stable && b1_prev);
    wire b1_holding = b1_stable;

    wire b2_pressed = (b2_stable && !b2_prev);
    wire b3_pressed = (b3_stable && !b3_prev);

    //==========================================================================
    // 7. ���� ���� (��ư0 + ��ư1 + ��ư2 + ��ư3)
    //==========================================================================
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            b0_prev <= 1'b0;
            b0_hold_counter <= 32'd0;
            b0_long_triggered <= 1'b0;
            btn1_held <= 1'b0;
            
            b1_prev <= 1'b0;
            b1_repeat_counter <= 32'd0;
            b1_first_dot_sent <= 1'b0;
            
            b2_prev <= 1'b0;
            b3_prev <= 1'b0;
            
            key_valid <= 1'b0;
            key_packet <= 11'd0;
            btn2_dot_pulse <= 1'b0;
        end else begin
            b0_prev <= b0_stable;
            b1_prev <= b1_stable;
            b2_prev <= b2_stable;
            b3_prev <= b3_stable;
            
            // �⺻��
            key_valid <= 1'b0;
            btn2_dot_pulse <= 1'b0;
            
            // ========== btn[2] ó�� (PAUSE) ==========
            if(b2_pressed) begin
                key_valid <= 1'b1;
                key_packet <= {TYPE_KEY, KEY_PAUSE};
            end
            
            // ========== btn[3] ó�� (CLEAR) ==========
            if(b3_pressed) begin
                key_valid <= 1'b1;
                key_packet <= {TYPE_KEY, KEY_CLEAR};
            end
            
            // ========== ��ư2 ó�� (btn[1] - DOT �ڵ� �ݺ�) ==========
            if(b1_pressed) begin
                b1_repeat_counter <= 32'd0;
                b1_first_dot_sent <= 1'b1;
                
                key_valid <= 1'b1;
                key_packet <= {TYPE_KEY, KEY_DOT};
                btn2_dot_pulse <= 1'b1;
            end
            else if(b1_holding && b1_first_dot_sent) begin
                if(b1_repeat_counter >= DIT_GAP_CYCLES) begin
                    b1_repeat_counter <= 32'd0;
                    
                    key_valid <= 1'b1;
                    key_packet <= {TYPE_KEY, KEY_DOT};
                    btn2_dot_pulse <= 1'b1;
                end else begin
                    b1_repeat_counter <= b1_repeat_counter + 1;
                end
            end
            else if(b1_released) begin
                b1_repeat_counter <= 32'd0;
                b1_first_dot_sent <= 1'b0;
            end
            
            // ========== ��ư1 ó�� (btn[0] - DOT/DASH) ==========
            if(b0_pressed) begin
                btn1_held <= 1'b1;
                b0_hold_counter <= 32'd0;
                b0_long_triggered <= 1'b0;
            end
            else if(b0_holding) begin
                if(!b0_long_triggered) begin
                    if(b0_hold_counter >= LONG_KEY_CYCLES) begin
                        b0_long_triggered <= 1'b1;
                        btn1_held <= 1'b0;
                        
                        key_valid <= 1'b1;
                        key_packet <= {TYPE_KEY, KEY_DASH};
                    end else begin
                        b0_hold_counter <= b0_hold_counter + 1;
                    end
                end
            end
            else if(b0_released) begin
                btn1_held <= 1'b0;
                
                if(!b0_long_triggered) begin
                    key_valid <= 1'b1;
                    key_packet <= {TYPE_KEY, KEY_DOT};
                end
                
                b0_hold_counter <= 32'd0;
                b0_long_triggered <= 1'b0;
            end
        end
    end

endmodule

//==========================================================================
// PiezoToneController - �ǿ��� ��Ʈ�ѷ� (���� ����)
//==========================================================================
module PiezoToneController (
    input  wire        clk,
    input  wire        rst_n,
    input  wire        btn1_held,                  // ��ư1 ������ ��
    input  wire        btn2_dot_pulse,             // ��ư2 DOT �޽�
    
    input  wire [31:0] dash_cycles,                // ��� �� ��
    input  wire [31:0] autorepeat_cycles,          // ��� �� ��
    
    input  wire        char_complete_beep,         // ���� �Ϸ� ������
    
    output reg         piezo_out
);

    parameter CLK_HZ = 25_000_000;
    
    // 440Hz �� (��ư1 ������ ��, ��ư2 DOT)
    parameter TONE_440HZ = 440;
    localparam TOGGLE_COUNT_440 = CLK_HZ / (2 * TONE_440HZ);
    
    // 220Hz �� (���� �Ϸ�)
    parameter TONE_220HZ = 220;
    localparam TOGGLE_COUNT_220 = CLK_HZ / (2 * TONE_220HZ);
    
    // ������ ���� �ð�
    localparam CHAR_BEEP_DURATION = CLK_HZ / 10;      // 100ms (���� �Ϸ�)
    localparam DOT_BEEP_DURATION = CLK_HZ / 20;       // 50ms (��ư2 DOT)
    
    reg [31:0] tone_counter;
    reg        tone_toggle;
    
    reg        char_beep_active;
    reg [31:0] char_beep_counter;
    
    reg        dot_beep_active;
    reg [31:0] dot_beep_counter;
    
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            tone_counter <= 32'd0;
            tone_toggle <= 1'b0;
            piezo_out <= 1'b0;
            char_beep_active <= 1'b0;
            char_beep_counter <= 32'd0;
            dot_beep_active <= 1'b0;
            dot_beep_counter <= 32'd0;
        end
        else begin
            // ���� �Ϸ� ������ Ʈ���� (�ֿ켱)
            if(char_complete_beep) begin
                char_beep_active <= 1'b1;
                char_beep_counter <= 32'd0;
                dot_beep_active <= 1'b0;      // �� �߰�
                dot_beep_counter <= 32'd0;    // �� �߰�
                tone_counter <= 32'd0;
                tone_toggle <= 1'b0;
            end
            // ��ư2 DOT ������ Ʈ����
            else if(btn2_dot_pulse) begin     // �� if �� else if ����
                dot_beep_active <= 1'b1;
                dot_beep_counter <= 32'd0;
                tone_counter <= 32'd0;
                tone_toggle <= 1'b0;
            end
            
            // �켱����: ���� �Ϸ� ������ > ��ư2 DOT ������ > ��ư1 ������
            if(char_beep_active) begin
                // ���� �Ϸ� ������ (220Hz, 100ms)
                if(char_beep_counter < CHAR_BEEP_DURATION) begin
                    char_beep_counter <= char_beep_counter + 1;
                    
                    if(tone_counter < TOGGLE_COUNT_220) begin
                        tone_counter <= tone_counter + 1;
                    end
                    else begin
                        tone_counter <= 32'd0;
                        tone_toggle <= ~tone_toggle;
                    end
                    piezo_out <= tone_toggle;
                end
                else begin
                    char_beep_active <= 1'b0;
                    piezo_out <= 1'b0;
                    tone_counter <= 32'd0;
                    tone_toggle <= 1'b0;
                end
            end
            else if(dot_beep_active) begin
                // ��ư2 DOT ������ (440Hz, 50ms)
                if(dot_beep_counter < DOT_BEEP_DURATION) begin
                    dot_beep_counter <= dot_beep_counter + 1;
                    
                    if(tone_counter < TOGGLE_COUNT_440) begin
                        tone_counter <= tone_counter + 1;
                    end
                    else begin
                        tone_counter <= 32'd0;
                        tone_toggle <= ~tone_toggle;
                    end
                    piezo_out <= tone_toggle;
                end
                else begin
                    dot_beep_active <= 1'b0;
                    piezo_out <= 1'b0;
                    tone_counter <= 32'd0;
                    tone_toggle <= 1'b0;
                end
            end
            else if(btn1_held) begin
                // ��ư1 ������ (440Hz)
                if(tone_counter < TOGGLE_COUNT_440) begin
                    tone_counter <= tone_counter + 1;
                end
                else begin
                    tone_counter <= 32'd0;
                    tone_toggle <= ~tone_toggle;
                end
                piezo_out <= tone_toggle;
            end
            else begin
                tone_counter <= 32'd0;
                tone_toggle <= 1'b0;
                piezo_out <= 1'b0;
            end
        end
    end

endmodule

module ServoController #(
    parameter CLK_HZ = 25_000_000
)(
    input  wire       clk,
    input  wire       rst_n,
    input  wire [8:0] angle,      // 0~180��
    output reg        pwm_out
);

    // PWM �ֱ�: 20ms (50Hz)
    localparam PWM_PERIOD = CLK_HZ / 50;  // 2,000,000 cycles
    
    // �޽� ��: 1ms(0��) ~ 2ms(180��) - ǥ�� ����
    localparam MIN_PULSE = CLK_HZ / 1000;  // 1ms = 100,000 cycles
    localparam MAX_PULSE = CLK_HZ / 500;   // 2ms = 200,000 cycles
    localparam PULSE_RANGE = MAX_PULSE - MIN_PULSE;  // 100,000 cycles
    
    reg [31:0] counter;
    reg [31:0] pulse_width;
    
    // ���� �� �޽� �� ��ȯ (�����Ҽ��� ����)
    // pulse_width = MIN_PULSE + (angle * PULSE_RANGE / 180)
    always @(*) begin
        // ���е� ���: (angle * PULSE_RANGE) ���� ���
        pulse_width = MIN_PULSE + ((angle * PULSE_RANGE) / 180);
    end
    
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            counter <= 32'd0;
            pwm_out <= 1'b0;
        end
        else begin
            if(counter < PWM_PERIOD - 1) begin
                counter <= counter + 1;
            end
            else begin
                counter <= 32'd0;
            end
            
            // PWM ���
            pwm_out <= (counter < pulse_width) ? 1'b1 : 1'b0;
        end
    end

endmodule

`timescale 1ns / 1ps

//==============================================================================
// LCD_Controller.v
// 16x2 Character LCD ���� ��� (HD44780 ȣȯ)
//==============================================================================
// ���:
// - DecodeUI�κ��� ���� ��� ��û ����
// - LCD �ʱ�ȭ �� ���� ���
// - 4��Ʈ ��� ����
//==============================================================================

`timescale 1ns / 1ps

module LCD_Controller #(
    parameter integer CLK_HZ = 25_000_000
)(
    input  wire        clk,
    input  wire        rst_n,
    
    // DecodeUI �������̽�
    input  wire        lcd_req,
    input  wire [1:0]  lcd_row,
    input  wire [3:0]  lcd_col,
    input  wire [7:0]  lcd_char,
    
    output reg         lcd_busy,
    output reg         lcd_done,
    
    // LCD �ϵ���� �� (8��Ʈ ���)
    output reg         lcd_e,
    output reg         lcd_rs,
    output reg         lcd_rw,
    output reg  [7:0]  lcd_data
);

    //==========================================================================
    // Ÿ�̹� ��� (CLK_HZ ����)
    //==========================================================================
    localparam integer CNT_15MS  = (CLK_HZ / 1000) * 15;      // 15ms
    localparam integer CNT_5MS   = (CLK_HZ / 1000) * 5;       // 5ms
    localparam integer CNT_100US = (CLK_HZ / 1_000_000) * 100; // 100us
    localparam integer CNT_CMD   = (CLK_HZ / 1_000_000) * 50;  // 50us
    localparam integer CNT_CLR   = (CLK_HZ / 1000) * 2;       // 2ms
    
    localparam integer E_PULSE_START = 2;
    localparam integer E_PULSE_END   = 22;
    localparam integer E_PULSE_TOTAL = E_PULSE_END + CNT_CMD;

    //==========================================================================
    // ��ɾ� ����
    //==========================================================================
    localparam [7:0] CMD_WAKEUP     = 8'h30;
    localparam [7:0] CMD_FUNC_SET   = 8'h38; // 8-bit, 2-line, 5x8 font
    localparam [7:0] CMD_DISP_OFF   = 8'h08;
    localparam [7:0] CMD_DISP_CLEAR = 8'h01;
    localparam [7:0] CMD_ENTRY_MODE = 8'h06; // Auto Increment
    localparam [7:0] CMD_DISP_ON    = 8'h0C; // Display On, Cursor Off

    //==========================================================================
    // ���� �ӽ�
    //==========================================================================
    localparam [4:0] ST_PWR_WAIT   = 0;
    localparam [4:0] ST_INIT_1     = 1;
    localparam [4:0] ST_INIT_2     = 2;
    localparam [4:0] ST_INIT_3     = 3;
    localparam [4:0] ST_FUNC_SET   = 4;
    localparam [4:0] ST_DISP_OFF   = 5;
    localparam [4:0] ST_DISP_CLR   = 6;
    localparam [4:0] ST_ENTRY_MODE = 7;
    localparam [4:0] ST_DISP_ON    = 8;
    localparam [4:0] ST_IDLE       = 9;
    localparam [4:0] ST_SET_ADDR   = 10;
    localparam [4:0] ST_WRITE_CHAR = 11;

    reg [4:0]  state;
    reg [31:0] wait_cnt;
    reg [6:0]  target_addr;

    //==========================================================================
    // �ʱ�ȭ �� ���� �ӽ�
    //==========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= ST_PWR_WAIT;
            wait_cnt <= 0;
            lcd_e <= 0;
            lcd_rs <= 0;
            lcd_rw <= 0;
            lcd_data <= 0;
            lcd_busy <= 1;
            lcd_done <= 0;
            target_addr <= 0;
        end else begin
            // �⺻��
            lcd_done <= 0;
            
            case (state)
                //==============================================================
                // �ʱ�ȭ ������ (����� �ڵ� ��Ÿ��)
                //==============================================================
                ST_PWR_WAIT: begin
                    lcd_busy <= 1;
                    if (wait_cnt >= CNT_15MS) begin
                        wait_cnt <= 0;
                        state <= ST_INIT_1;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_INIT_1: begin // 0x30
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_WAKEUP;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= (CNT_5MS + E_PULSE_END)) begin
                        wait_cnt <= 0;
                        state <= ST_INIT_2;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_INIT_2: begin // 0x30
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_WAKEUP;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= (CNT_100US + E_PULSE_END)) begin
                        wait_cnt <= 0;
                        state <= ST_INIT_3;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_INIT_3: begin // 0x30
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_WAKEUP;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        state <= ST_FUNC_SET;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_FUNC_SET: begin // 0x38
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_FUNC_SET;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        state <= ST_DISP_OFF;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_DISP_OFF: begin // 0x08
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_DISP_OFF;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        state <= ST_DISP_CLR;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_DISP_CLR: begin // 0x01
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_DISP_CLEAR;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= (CNT_CLR + E_PULSE_END)) begin
                        wait_cnt <= 0;
                        state <= ST_ENTRY_MODE;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_ENTRY_MODE: begin // 0x06
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_ENTRY_MODE;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        state <= ST_DISP_ON;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_DISP_ON: begin // 0x0C
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= CMD_DISP_ON;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        lcd_busy <= 0;
                        state <= ST_IDLE;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                //==============================================================
                // ��� �� ���� ���
                //==============================================================
                ST_IDLE: begin
                    lcd_e <= 0;
                    lcd_busy <= 0;
                    wait_cnt <= 0;
                    
                    if (lcd_req) begin
                        lcd_busy <= 1;
                        
                        // ��ǥ ���
                        if (lcd_row == 2'b00) begin
                            target_addr <= {3'b000, lcd_col}; // 0x00 + col
                        end else begin
                            target_addr <= {3'b100, lcd_col}; // 0x40 + col
                        end
                        
                        state <= ST_SET_ADDR;
                    end
                end

                ST_SET_ADDR: begin
                    lcd_rs <= 0;
                    lcd_rw <= 0;
                    lcd_data <= {1'b1, target_addr}; // 0x80 | Address
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        state <= ST_WRITE_CHAR;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                ST_WRITE_CHAR: begin
                    lcd_rs <= 1; // Data ���
                    lcd_rw <= 0;
                    lcd_data <= lcd_char;
                    
                    if (wait_cnt == E_PULSE_START) lcd_e <= 1;
                    else if (wait_cnt == E_PULSE_END) lcd_e <= 0;
                    
                    if (wait_cnt >= E_PULSE_TOTAL) begin
                        wait_cnt <= 0;
                        lcd_done <= 1;
                        lcd_busy <= 0;
                        state <= ST_IDLE;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end

                default: state <= ST_PWR_WAIT;
            endcase
        end
    end

endmodule