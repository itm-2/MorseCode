//==============================================================================
// Piezo Controller Module (PWM Generator)
//==============================================================================
module piezo_controller (
    input wire clk,              // 50MHz
    input wire rst_n,
    
    // Control Interface
    input wire enable,           // Piezo Ȱ��ȭ
    input wire [15:0] duration,  // ���� �ð� (ms ����)
    input wire [15:0] frequency, // ���ļ� (Hz ����)
    
    // PWM Output
    output reg pwm_out
);

//==============================================================================
// Parameters
//==============================================================================
localparam CLK_FREQ = 50_000_000;  // 50MHz

//==============================================================================
// Internal Registers
//==============================================================================
reg [31:0] duration_counter;   // ���� �ð� ī���� (Ŭ�� ����Ŭ)
reg [31:0] period_counter;     // PWM �ֱ� ī����
reg [31:0] half_period;        // ���ֱ� (Ŭ�� ����Ŭ)
reg [31:0] total_duration;     // �� ���� �ð� (Ŭ�� ����Ŭ)
reg active;                    // ���� Ȱ�� ����

//==============================================================================
// Duration & Period Calculation
//==============================================================================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        half_period <= 32'd25000;      // �⺻��: 1kHz (50MHz / 2000)
        total_duration <= 32'd50000;   // �⺻��: 1ms
    end else if (enable && !active) begin
        // ���ֱ� ���: CLK_FREQ / (2 * frequency)
        half_period <= CLK_FREQ / (frequency << 1);
        
        // �� ���� �ð� ���: duration(ms) * CLK_FREQ / 1000
        total_duration <= (duration * (CLK_FREQ / 1000));
    end
end

//==============================================================================
// PWM Generation Logic
//==============================================================================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        pwm_out <= 1'b0;
        duration_counter <= 32'b0;
        period_counter <= 32'b0;
        active <= 1'b0;
        
    end else begin
        if (enable && !active) begin
            // ���ο� �� ����
            active <= 1'b1;
            duration_counter <= 32'b0;
            period_counter <= 32'b0;
            pwm_out <= 1'b1;
            
        end else if (active) begin
            // ���� �ð� üũ
            if (duration_counter >= total_duration) begin
                // ���� �ð� ����
                active <= 1'b0;
                pwm_out <= 1'b0;
                duration_counter <= 32'b0;
                period_counter <= 32'b0;
                
            end else begin
                // PWM ���
                if (period_counter >= half_period) begin
                    pwm_out <= ~pwm_out;
                    period_counter <= 32'b0;
                end else begin
                    period_counter <= period_counter + 1;
                end
                
                duration_counter <= duration_counter + 1;
            end
        end else begin
            pwm_out <= 1'b0;
        end
    end
end

endmodule