`timescale 1ns / 1ps

module Button_Debouncer (
    input wire clk,       // [�ý��� ǥ��] 100kHz Ŭ�� �Է�
    input wire rst_n,     // Active Low Reset
    input wire btn_in,    // ����� ���� ��ư �Է�
    output reg btn_out    // ��ٿ�� �Ϸ�� ������ ���
);

    // =========================================================================
    // 1. �Ķ���� ���� (100kHz ����)
    // =========================================================================
    parameter CLK_FREQ    = 100_000; // 100kHz
    parameter DEBOUNCE_MS = 20;      // 20ms
    
    // ��ǥ ī��Ʈ: 100,000 * 0.02 = 2,000
    localparam CNT_MAX = (CLK_FREQ / 1000) * DEBOUNCE_MS;

    // =========================================================================
    // 2. ���� ����
    // =========================================================================
    reg [31:0] cnt;
    reg btn_sync_0;       // ��ũ�γ����� 1
    reg btn_sync_1;       // ��ũ�γ����� 2

    // =========================================================================
    // 3. ���� ����
    // =========================================================================
    
    // 3-1. �Է� ����ȭ (�ܺ� ��ȣ -> ���� Ŭ��)
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            btn_sync_0 <= 1'b0;
            btn_sync_1 <= 1'b0;
        end else begin
            btn_sync_0 <= btn_in;
            btn_sync_1 <= btn_sync_0;
        end
    end

    // 3-2. ��ٿ�� ī����
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cnt <= 0;
            btn_out <= 1'b0;
        end else begin
            // ���� ��°� �Է�(����ȭ��)�� �ٸ��� ī��Ʈ ����
            if (btn_out != btn_sync_1) begin
                cnt <= cnt + 1;
                
                // 20ms(2000Ŭ��) ���� �����Ǹ� �� ����
                if (cnt >= CNT_MAX) begin
                    btn_out <= btn_sync_1;
                    cnt <= 0;
                end
            end else begin
                // �߰��� ���� Ƣ�� ī���� �ʱ�ȭ
                cnt <= 0;
            end
        end
    end

endmodule